`include "i2s.v"
//NOTES:

module peddle(data_in, data_out);

//need an i2s_rx(data_in)

//need clk_div module

//need pwm(data_out)

//need buffers



endmodule

module pwm();

endmodule
